magic
tech sky130A
timestamp 1633032407
<< error_p >>
rect -535 1149 -518 1150
rect -535 1130 -518 1131
rect -104 -37 -87 -36
rect 134 -39 151 -38
rect 21 -407 38 -406
<< nwell >>
rect -2673 6125 2341 7034
rect -185 200 86 6125
rect -286 -136 347 200
<< pwell >>
rect -1557 194 -1031 320
<< nmos >>
rect -1344 207 -1244 307
<< pmos >>
rect -27 -97 73 3
<< ndiff >>
rect -1544 281 -1344 307
rect -1544 229 -1535 281
rect -1483 229 -1344 281
rect -1544 207 -1344 229
rect -1244 279 -1044 307
rect -1244 228 -1117 279
rect -1065 228 -1044 279
rect -1244 207 -1044 228
<< pdiff >>
rect -123 -19 -27 3
rect -123 -37 -104 -19
rect -87 -37 -27 -19
rect -123 -53 -27 -37
rect -123 -71 -104 -53
rect -87 -71 -27 -53
rect -123 -97 -27 -71
rect 73 -21 177 3
rect 73 -39 134 -21
rect 151 -39 177 -21
rect 73 -55 177 -39
rect 73 -73 134 -55
rect 151 -73 177 -55
rect 73 -97 177 -73
<< ndiffc >>
rect -1535 229 -1483 281
rect -1117 228 -1065 279
<< pdiffc >>
rect -104 -37 -87 -19
rect -104 -71 -87 -53
rect 134 -39 151 -21
rect 134 -73 151 -55
<< nsubdiff >>
rect -545 6538 832 6592
rect -545 6419 -149 6538
rect 38 6419 832 6538
rect -545 6321 832 6419
<< nsubdiffcont >>
rect -149 6419 38 6538
<< poly >>
rect -1344 307 -1244 385
rect -1344 -43 -1244 207
rect -27 3 73 42
rect -1344 -60 -1301 -43
rect -1283 -60 -1244 -43
rect -1344 -115 -1244 -60
rect -27 -389 73 -97
rect -27 -407 21 -389
rect 38 -407 73 -389
rect -27 -423 73 -407
rect -27 -441 21 -423
rect 38 -441 73 -423
rect -27 -458 73 -441
<< polycont >>
rect -1301 -60 -1283 -43
rect 21 -407 38 -389
rect 21 -441 38 -423
<< xpolycontact >>
rect -1153 5717 -973 6081
rect -2355 4764 -2160 5124
rect 1178 5065 1341 5421
rect -1175 383 -995 747
rect 2039 4956 2208 5310
rect -2355 -482 -2160 -122
rect 1171 -163 1356 207
rect 2017 -496 2186 -142
<< xpolyres >>
rect -2306 -122 -2271 4764
rect -1092 747 -1057 5717
rect 1261 207 1296 5065
rect 2122 -142 2157 4956
<< locali >>
rect -2086 6666 1949 6737
rect -2086 6360 -1965 6666
rect -1588 6663 1949 6666
rect -1588 6538 1498 6663
rect -1588 6419 -149 6538
rect 38 6419 1498 6538
rect -1588 6360 1498 6419
rect -2086 6357 1498 6360
rect 1839 6357 1949 6663
rect -2086 6295 1949 6357
rect -1157 6081 -968 6295
rect -1157 6067 -1153 6081
rect -1159 5868 -1153 6067
rect -2711 5822 -1486 5828
rect -3412 5647 -1486 5822
rect -973 6067 -968 6081
rect -973 5868 -966 6067
rect -3412 5378 -3299 5647
rect -2994 5628 -1486 5647
rect -2994 5378 -1897 5628
rect -3412 5359 -1897 5378
rect -1592 5359 -1486 5628
rect 1614 5462 1880 6295
rect -3412 5222 -1486 5359
rect 671 5264 933 5276
rect -3412 5216 -2187 5222
rect -2364 5124 -2187 5216
rect 671 5151 1178 5264
rect -2364 4925 -2355 5124
rect -2160 4917 -1542 4943
rect -2160 4764 -1478 4917
rect -2344 4752 -1478 4764
rect -1657 281 -1478 4752
rect -598 1167 -450 1217
rect -598 1149 -535 1167
rect -518 1149 -450 1167
rect -598 1131 -450 1149
rect -598 1113 -535 1131
rect -518 1113 -450 1131
rect -598 655 -450 1113
rect 671 655 933 5151
rect 1614 5329 2183 5462
rect 1614 5317 1880 5329
rect 2031 5310 2176 5329
rect 2031 5127 2039 5310
rect -830 513 945 655
rect -1657 229 -1535 281
rect -1483 229 -1478 281
rect -1657 168 -1478 229
rect -1141 279 -1037 383
rect -1141 228 -1117 279
rect -1065 228 -1037 279
rect -1141 211 -1037 228
rect -1141 177 -1040 211
rect -1321 9 -68 10
rect -1365 2 -68 9
rect 108 2 1171 12
rect -1365 -19 -55 2
rect -1365 -37 -104 -19
rect -87 -37 -55 -19
rect -1365 -43 -55 -37
rect -1365 -60 -1301 -43
rect -1283 -53 -55 -43
rect -1283 -60 -104 -53
rect -1365 -71 -104 -60
rect -87 -71 -55 -53
rect -1365 -97 -55 -71
rect 107 -21 1171 2
rect 107 -39 134 -21
rect 151 -39 1171 -21
rect 107 -55 1171 -39
rect 107 -73 134 -55
rect 151 -73 1171 -55
rect 107 -97 1171 -73
rect -1365 -99 -68 -97
rect 108 -109 1171 -97
rect -2466 -454 -2355 -360
rect -2160 -365 -2138 -360
rect -2160 -368 33 -365
rect -2160 -389 2017 -368
rect -2160 -407 21 -389
rect 38 -407 2017 -389
rect -2160 -423 2017 -407
rect -2160 -441 21 -423
rect 38 -441 2017 -423
rect -2160 -451 2017 -441
rect -2160 -454 79 -451
rect -30 -754 79 -454
rect 2186 -451 2227 -368
rect -30 -772 3 -754
rect 20 -772 39 -754
rect 56 -772 79 -754
rect -30 -805 79 -772
<< viali >>
rect -1965 6360 -1588 6666
rect 1498 6357 1839 6663
rect -3299 5378 -2994 5647
rect -1897 5359 -1592 5628
rect -535 1149 -518 1167
rect -535 1113 -518 1131
rect 3 -772 20 -754
rect 39 -772 56 -754
<< metal1 >>
rect -2086 6666 1949 6737
rect -2086 6360 -1965 6666
rect -1588 6663 1949 6666
rect -1588 6360 1498 6663
rect -2086 6357 1498 6360
rect 1839 6357 1949 6663
rect -2086 6295 1949 6357
rect -2711 5822 -1486 5828
rect -3412 5647 -1486 5822
rect -3412 5378 -3299 5647
rect -2994 5628 -1486 5647
rect -2994 5378 -1897 5628
rect -3412 5359 -1897 5378
rect -1592 5359 -1486 5628
rect -3412 5222 -1486 5359
rect -3412 5216 -2187 5222
rect -598 1167 -462 1211
rect -598 1149 -535 1167
rect -518 1149 -462 1167
rect -598 1131 -462 1149
rect -598 1113 -535 1131
rect -518 1113 -462 1131
rect -598 1075 -462 1113
rect -50 -754 109 -714
rect -50 -772 3 -754
rect 20 -772 39 -754
rect 56 -772 109 -754
rect -50 -811 109 -772
<< labels >>
rlabel metal1 s 3 -786 58 -740 4 vin
port 1 nsew
rlabel metal1 s -548 1112 -505 1168 4 vout
port 2 nsew
rlabel metal1 s -255 6390 143 6617 4 vdd
port 3 nsew
rlabel metal1 s -2648 5354 -2269 5582 4 gnd
port 4 nsew
<< end >>
